mquinto@hpmichele.dyndns.cern.ch.10823:1484041098