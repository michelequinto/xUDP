package test_pkg;
   
`include <uvm_macros.svh>

import uvm_pkg::*;
import mvc_pkg::*;
import mgc_ethernet_v1_0_pkg::*;
import env_pkg::*;

`include "ethernet_upper_layer_packet_seq.svh"
`include "ethernet_monitors.svh"

endpackage
